`timescale 1ns/1ps
// Bus interface unit: assumes two branches of the bus -
// 1. connect to dmem
// 2. connect to a single peripheral
// The BIU needs to know the addresses at which DMEM and peripheral are
// connected, so it can do the required multiplexing. 
// These need to be added as part of your code. 
module biu (
    input clk,
    input reset,
    input [31:0] daddr,
    input [31:0] dwdata,
    input [3:0] dwe,
    output [31:0] drdata,

    // Signals going to/from dmem
    output [31:0] daddr1,
    output [31:0] dwdata1,
    output [3:0]  dwe1,
    input  [31:0] drdata1,

    // Signals going to/from peripheral
    output [31:0] daddr2,
    output [31:0] dwdata2,
    output [3:0]  dwe2,
    input  [31:0] drdata2
);
    reg[31:0] daddr1,dwdata1,daddr2,dwdata2;
    reg[3:0] dwe1,dwe2;

    // Modify below so that depending on the actual daddr range the BIU decides whether 
    // the response was from DMEM or peripheral - maybe a MUX?
    assign drdata = drdata1;

    // Send values to DMEM or peripheral (or both if it does not matter)
    // as required    

//     initial begin
//         if (daddr == 0x34560)
//             $monitor($time);
//     end
    
    always@(*)
        begin
    
            if (daddr == 32'h00034560)
                begin
//                    $display("Inside perifh");
                    daddr2 = daddr;
                    dwdata2 = dwdata;
                    dwe2 = dwe;
                end
            else
                begin
                    //$display("Inside dmem");                    
                    daddr1 = daddr;
                    dwdata1 = dwdata;
                    dwe1 = dwe;
                end
        end
    
endmodule